module top_module ( input a, input b, output out );
    mod_a instance1 (a, b, out); 
    //É como declarar uma função em c só que em verilog;
endmodule
